`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:	-
// Engineer: Ahmet Alparslan Celik
// 
// Create Date:    22:25:41 12/12/2015  
// Design Name: 	-
// Module Name:    rom_glcd 
// Project Name: 	FPGA implementation of simple XOR cipher
// Target Devices: -
// Tool versions: -
// Description: -
//
// Dependencies: -
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module rom_glcd
	(
		input clk, reset,
		input [6:0] R_A,
		output [39:0] R_D 
	);
	
	reg [39:0] ROM [95:0];
	
	assign R_D = ROM[R_A];
	
	always@(posedge clk)
		if(reset==1'b0) 
			begin
				ROM[0] <= {8'h00, 8'h00, 8'h00, 8'h00, 8'h00}; // 20  
				ROM[1] <= {8'h00, 8'h00, 8'h5f, 8'h00, 8'h00}; // 21 !
				ROM[2] <= {8'h00, 8'h07, 8'h00, 8'h07, 8'h00}; // 22 "
				ROM[3] <= {8'h14, 8'h7f, 8'h14, 8'h7f, 8'h14}; // 23 #
				ROM[4] <= {8'h24, 8'h2a, 8'h7f, 8'h2a, 8'h12}; // 24 $
				ROM[5] <= {8'h23, 8'h13, 8'h08, 8'h64, 8'h62}; // 25 %
				ROM[6] <= {8'h36, 8'h49, 8'h55, 8'h22, 8'h50}; // 26 &
				ROM[7] <= {8'h00, 8'h05, 8'h03, 8'h00, 8'h00}; // 27 '
				ROM[8] <= {8'h00, 8'h1c, 8'h22, 8'h41, 8'h00}; // 28 (
				ROM[9] <= {8'h00, 8'h41, 8'h22, 8'h1c, 8'h00}; // 29 )
				ROM[10] <= {8'h14, 8'h08, 8'h3e, 8'h08, 8'h14}; // 2a *
				ROM[11] <= {8'h08, 8'h08, 8'h3e, 8'h08, 8'h08}; // 2b +
				ROM[12] <= {8'h00, 8'h50, 8'h30, 8'h00, 8'h00}; // 2c ,
				ROM[13] <= {8'h08, 8'h08, 8'h08, 8'h08, 8'h08}; // 2d -
				ROM[14] <= {8'h00, 8'h60, 8'h60, 8'h00, 8'h00}; // 2e .
				ROM[15] <= {8'h20, 8'h10, 8'h08, 8'h04, 8'h02}; // 2f /
				ROM[16] <= {8'h3e, 8'h51, 8'h49, 8'h45, 8'h3e}; // 30 0
				ROM[17] <= {8'h00, 8'h42, 8'h7f, 8'h40, 8'h00}; // 31 1
				ROM[18] <= {8'h42, 8'h61, 8'h51, 8'h49, 8'h46}; // 32 2
				ROM[19] <= {8'h21, 8'h41, 8'h45, 8'h4b, 8'h31}; // 33 3
				ROM[20] <= {8'h18, 8'h14, 8'h12, 8'h7f, 8'h10}; // 34 4
				ROM[21] <= {8'h27, 8'h45, 8'h45, 8'h45, 8'h39}; // 35 5
				ROM[22] <= {8'h3c, 8'h4a, 8'h49, 8'h49, 8'h30}; // 36 6
				ROM[23] <= {8'h01, 8'h71, 8'h09, 8'h05, 8'h03}; // 37 7
				ROM[24] <= {8'h36, 8'h49, 8'h49, 8'h49, 8'h36}; // 38 8
				ROM[25] <= {8'h06, 8'h49, 8'h49, 8'h29, 8'h1e}; // 39 9
				ROM[26] <= {8'h00, 8'h36, 8'h36, 8'h00, 8'h00}; // 3a :
				ROM[27] <= {8'h00, 8'h56, 8'h36, 8'h00, 8'h00}; // 3b ;
				ROM[28] <= {8'h08, 8'h14, 8'h22, 8'h41, 8'h00}; // 3c <
				ROM[29] <= {8'h14, 8'h14, 8'h14, 8'h14, 8'h14}; // 3d =
				ROM[30] <= {8'h00, 8'h41, 8'h22, 8'h14, 8'h08}; // 3e >
				ROM[31] <= {8'h02, 8'h01, 8'h51, 8'h09, 8'h06}; // 3f ?
				ROM[32] <= {8'h32, 8'h49, 8'h79, 8'h41, 8'h3e}; // 40 @
				ROM[33] <= {8'h7e, 8'h11, 8'h11, 8'h11, 8'h7e}; // 41 A
				ROM[34] <= {8'h7f, 8'h49, 8'h49, 8'h49, 8'h36}; // 42 B
				ROM[35] <= {8'h3e, 8'h41, 8'h41, 8'h41, 8'h22}; // 43 C
				ROM[36] <= {8'h7f, 8'h41, 8'h41, 8'h22, 8'h1c}; // 44 D
				ROM[37] <= {8'h7f, 8'h49, 8'h49, 8'h49, 8'h41}; // 45 E
				ROM[38] <= {8'h7f, 8'h09, 8'h09, 8'h09, 8'h01}; // 46 F
				ROM[39] <= {8'h3e, 8'h41, 8'h49, 8'h49, 8'h7a}; // 47 G
				ROM[40] <= {8'h7f, 8'h08, 8'h08, 8'h08, 8'h7f}; // 48 H
				ROM[41] <= {8'h00, 8'h41, 8'h7f, 8'h41, 8'h00}; // 49 I
				ROM[42] <= {8'h20, 8'h40, 8'h41, 8'h3f, 8'h01}; // 4a J
				ROM[43] <= {8'h7f, 8'h08, 8'h14, 8'h22, 8'h41}; // 4b K
				ROM[44] <= {8'h7f, 8'h40, 8'h40, 8'h40, 8'h40}; // 4c L
				ROM[45] <= {8'h7f, 8'h02, 8'h0c, 8'h02, 8'h7f}; // 4d M
				ROM[46] <= {8'h7f, 8'h04, 8'h08, 8'h10, 8'h7f}; // 4e N
				ROM[47] <= {8'h3e, 8'h41, 8'h41, 8'h41, 8'h3e}; // 4f O
				ROM[48] <= {8'h7f, 8'h09, 8'h09, 8'h09, 8'h06}; // 50 P
				ROM[49] <= {8'h3e, 8'h41, 8'h51, 8'h21, 8'h5e}; // 51 Q
				ROM[50] <= {8'h7f, 8'h09, 8'h19, 8'h29, 8'h46}; // 52 R
				ROM[51] <= {8'h46, 8'h49, 8'h49, 8'h49, 8'h31}; // 53 S
				ROM[52] <= {8'h01, 8'h01, 8'h7f, 8'h01, 8'h01}; // 54 T
				ROM[53] <= {8'h3f, 8'h40, 8'h40, 8'h40, 8'h3f}; // 55 U
				ROM[54] <= {8'h1f, 8'h20, 8'h40, 8'h20, 8'h1f}; // 56 V
				ROM[55] <= {8'h3f, 8'h40, 8'h38, 8'h40, 8'h3f}; // 57 W
				ROM[56] <= {8'h63, 8'h14, 8'h08, 8'h14, 8'h63}; // 58 X
				ROM[57] <= {8'h07, 8'h08, 8'h70, 8'h08, 8'h07}; // 59 Y
				ROM[58] <= {8'h61, 8'h51, 8'h49, 8'h45, 8'h43}; // 5a Z
				ROM[59] <= {8'h00, 8'h7f, 8'h41, 8'h41, 8'h00}; // 5b [
				ROM[60] <= {8'h02, 8'h04, 8'h08, 8'h10, 8'h20}; // 5c \
				ROM[61] <= {8'h00, 8'h41, 8'h41, 8'h7f, 8'h00}; // 5d ]
				ROM[62] <= {8'h04, 8'h02, 8'h01, 8'h02, 8'h04}; // 5e ^
				ROM[63] <= {8'h40, 8'h40, 8'h40, 8'h40, 8'h40}; // 5f _
				ROM[64] <= {8'h00, 8'h01, 8'h02, 8'h04, 8'h00}; // 60 `
				ROM[65] <= {8'h20, 8'h54, 8'h54, 8'h54, 8'h78}; // 61 a
				ROM[66] <= {8'h7f, 8'h48, 8'h44, 8'h44, 8'h38}; // 62 b
				ROM[67] <= {8'h38, 8'h44, 8'h44, 8'h44, 8'h20}; // 63 c
				ROM[68] <= {8'h38, 8'h44, 8'h44, 8'h48, 8'h7f}; // 64 d
				ROM[69] <= {8'h38, 8'h54, 8'h54, 8'h54, 8'h18}; // 65 e
				ROM[70] <= {8'h08, 8'h7e, 8'h09, 8'h01, 8'h02}; // 66 f
				ROM[71] <= {8'h0c, 8'h52, 8'h52, 8'h52, 8'h3e}; // 67 g
				ROM[72] <= {8'h7f, 8'h08, 8'h04, 8'h04, 8'h78}; // 68 h
				ROM[73] <= {8'h00, 8'h44, 8'h7d, 8'h40, 8'h00}; // 69 i
				ROM[74] <= {8'h20, 8'h40, 8'h44, 8'h3d, 8'h00}; // 6a j 
				ROM[75] <= {8'h7f, 8'h10, 8'h28, 8'h44, 8'h00}; // 6b k
				ROM[76] <= {8'h00, 8'h41, 8'h7f, 8'h40, 8'h00}; // 6c l
				ROM[77] <= {8'h7c, 8'h04, 8'h18, 8'h04, 8'h78}; // 6d m
				ROM[78] <= {8'h7c, 8'h08, 8'h04, 8'h04, 8'h78}; // 6e n
				ROM[79] <= {8'h38, 8'h44, 8'h44, 8'h44, 8'h38}; // 6f o
				ROM[80] <= {8'h7c, 8'h14, 8'h14, 8'h14, 8'h08}; // 70 p
				ROM[81] <= {8'h08, 8'h14, 8'h14, 8'h18, 8'h7c}; // 71 q
				ROM[82] <= {8'h7c, 8'h08, 8'h04, 8'h04, 8'h08}; // 72 r
				ROM[83] <= {8'h48, 8'h54, 8'h54, 8'h54, 8'h20}; // 73 s
				ROM[84] <= {8'h04, 8'h3f, 8'h44, 8'h40, 8'h20}; // 74 t
				ROM[85] <= {8'h3c, 8'h40, 8'h40, 8'h20, 8'h7c}; // 75 u
				ROM[86] <= {8'h1c, 8'h20, 8'h40, 8'h20, 8'h1c}; // 76 v
				ROM[87] <= {8'h3c, 8'h40, 8'h30, 8'h40, 8'h3c}; // 77 w
				ROM[88] <= {8'h44, 8'h28, 8'h10, 8'h28, 8'h44}; // 78 x
				ROM[89] <= {8'h0c, 8'h50, 8'h50, 8'h50, 8'h3c}; // 79 y
				ROM[90] <= {8'h44, 8'h64, 8'h54, 8'h4c, 8'h44}; // 7a z
				ROM[91] <= {8'h00, 8'h08, 8'h36, 8'h41, 8'h00}; // 7b {
				ROM[92] <= {8'h00, 8'h00, 8'h7f, 8'h00, 8'h00}; // 7c |
				ROM[93] <= {8'h00, 8'h41, 8'h36, 8'h08, 8'h00}; // 7d }
				ROM[94] <= {8'h10, 8'h08, 8'h08, 8'h10, 8'h08}; // 7e ~
				ROM[95] <= {8'h78, 8'h46, 8'h41, 8'h46, 8'h78}; // 7f DEL
			end
endmodule
